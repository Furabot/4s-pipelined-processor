`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 21.04.2020 18:59:51
// Design Name: 
// Module Name: processor_mc
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module processor_mc(
    input clk,
    input reset
    );
    
    wire [7:0] instruction_code_if; //instruction code from the IF stage
    wire [7:0] instruction_code; //instruction code from IF/ID register 
    wire [7:0] write_data; //write data from the WB stage
    wire [7:0] read_data1_id; 
    wire [7:0] read_data2_id; //register data from the register file
    wire regwrite; //regwrite control signal
    wire aluop_id; //aluop signal generated by the CU; input to ID/EX register
    wire shamt_sel_id; //shamt signal generated by the CU; input to ID/EX register
    wire regwrite_id; //regwrite signal generated by the CU; input to ID/EX register
    wire [7:0] shamt_id; //shift-amount, input into ID/EX register
    wire [7:0] regfile_data1; 
    wire [7:0] regfile_data2; //register file data 
    wire [7:0] shamt; //shift-amount
    wire aluop; //aluop control signal
    wire shamt_sel; //shamt control signal
    wire regwrite_ex; //regwrite singal, input to EX/WB register
    wire [2:0] prev_ins_dst_ex; //destination register, input to EX/WB register
    wire [2:0] curr_ins_s1; 
    wire [2:0] curr_ins_s2; //source registers
    wire [7:0] fwd_data; //data forwarded from WB stage
    wire fwdA; //control line to select the forwarded data for input 1 of ALU
    wire [7:0] alu_data1; //data input 1 to the ALU
    wire fwdB; //control line to select the forwarded data for input 2 of ALU
    wire [7:0] alu_data2; //data input 1 to the ALU
    wire [7:0] alu_result_ex; //ALU result, input to the EX/WB register
    wire alu_zero;
    wire [2:0] prev_ins_dst; //destination register
    
    assign shamt_id[7:3] = 5'b00000;
    assign shamt_id[2:0] = instruction_code[2:0]; //zero-padding shift-amount, to obtain 8-bit data
    assign fwd_data = write_data; //forwarded data = WB data
    
    //IF stage
    instruction_fetch IF(clk, reset, instruction_code_if); //instruction fetch unit
    IFID IFIDreg(clk, reset, instruction_code_if, instruction_code); //IF/ID register
    //ID stage
    register_file_noclk ID_regfile(instruction_code[5:3], instruction_code[2:0], prev_ins_dst, write_data, read_data1_id, read_data2_id, regwrite, reset); //register file                  
    control ID_cu(instruction_code[7:6], aluop_id, shamt_sel_id, regwrite_id); //control unit
    IDEX IDEXreg(clk, reset, read_data1_id, read_data2_id, shamt_id, aluop_id, shamt_sel_id, regwrite_id, instruction_code[5:3], instruction_code[5:3], instruction_code[2:0], regfile_data1, regfile_data2, shamt, aluop, shamt_sel, regwrite_ex, prev_ins_dst_ex, curr_ins_s1, curr_ins_s2); //IDEX register
    //EX,WB stage
    mux alu_mux1(regfile_data1, fwd_data, fwdA, alu_data1); //mux for input 1 of the ALU, to select register data or forwarded data
    mux3 alu_mux2(regfile_data2, fwd_data, shamt, shamt_sel, fwdB, alu_data2); //mux for input 2 of the ALU, to select register data, forwarded data or shift-amount data        
    alu alu(alu_data1, alu_data2, aluop, alu_result_ex, alu_zero); //ALU
    EXWB EXWBreg(clk, reset, alu_result_ex, regwrite_ex, prev_ins_dst_ex, write_data, regwrite, prev_ins_dst); //EX/WB register
    fwd forward_unit(prev_ins_dst, curr_ins_s1, curr_ins_s2, fwdA, fwdB); //forwarding unit
    
endmodule
